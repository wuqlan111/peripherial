
/****************************************************************************************
* Module Name:     spi_core
* Author:          wuqlan
* Email:           
* Date Created:    2023/4/2
* Description:     SPI core module.
*                  
*
* Version:         0.1
*****************************************************************************************/
module spi_core (

    /*-------system clk and reset signal*/
    input  clk_in,
    input  rstn_in,

    /*------spi signal------*/
    output   miso_out,
    input   miso_in,
    input  mosi_in,
    output  mosi_out,
    output  sck_in,
    input   sck_out,
    input  ss_in,
    output  ss_out

);











endmodule




