
/****************************************************************************************
* Module Name:     spi_top
* Author:          wuqlan
* Email:           
* Date Created:    2023/4/2
* Description:     SPI top module.
*                  
*
* Version:         0.1
*****************************************************************************************/
module   spi_top(

                input  clk_in,
                input  rstn_in,


                /*--------spi module top signal-------*/
                inout  miso_io,
                inout  mosi_in,
                inout  sck_in,
                inout  ss_io


                    );



















endmodule


